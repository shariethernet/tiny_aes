/*
 * Copyright 2012, Homer Hsing <homer.hsing@gmail.com>
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`timescale 1ns / 1ps

module test_aes_128;

	// Inputs
	reg clk;
	reg [127:0] state;
	reg [127:0] key;

	// Outputs
	wire [127:0] out;

	// Instantiate the Unit Under Test (UUT)
	aes_128 uut (
		.clk(clk), 
		.state(state), 
		.key(key), 
		.out(out)
	);

	initial begin
		clk = 0;
		state = 0;
		key = 0;
		#100;
        /*
         * TIMEGRP "key" OFFSET = IN 6.4 ns VALID 6 ns AFTER "clk" HIGH;
         * TIMEGRP "state" OFFSET = IN 6.4 ns VALID 6 ns AFTER "clk" HIGH;
         * TIMEGRP "out" OFFSET = OUT 2.2 ns BEFORE "clk" HIGH;
         */
        @ (negedge clk);
        # 2;
        state = 128'h3243f6a8_885a308d_313198a2_e0370734;
        key   = 128'h2b7e1516_28aed2a6_abf71588_09cf4f3c;
        #10;
        state = 128'h00112233_44556677_8899aabb_ccddeeff;
        key   = 128'h00010203_04050607_08090a0b_0c0d0e0f;
        #10;
        state = 128'h0;
        key   = 128'h0;
        #10;
        state = 128'h0;
        key   = 128'h1;
        #10;
        state = 128'h1;
        key   = 128'h0;
        #10;
 state = 128'h7369c667ec4aff51abbacd2946e3fbf2;
key =      128'hf854c27c8de7e81b632e5a769ac99f33;


#10;
 state = 128'hb70d32665aa3583117055d25d45ee958;
key =      128'hc6cdb2ab1154b49b4174820e87dc3d21;


#10;
 state = 128'ha13ee97067fce141977e013e966bdcea;
key =      128'h2a5c388ffb3bb0ec543caf325cdb18ec;


#10;
 state = 128'h43fe1a023aaafafbe6d129fb947c3c05;
key =      128'h61bed875bb5cf989950f99a8b3f1ebb1;


#10;
 state = 128'h00f7ef05e53aa1e9d0cb0bcabd644748;
key =      128'ha81e231fc5647b1cc55a731463794b5e;


#10;
 state = 128'h2464703bdc099e11f2acd4aa3baf101b;
key =      128'h50e3cd335c15474819226fbbf57d9bba;


#10;
 state = 128'h1c1ae10b29f8237f131ba4f8e84ecab5;
key =      128'he0383298343d4d79774e5fbc056ccbfa;


#10;
 state = 128'h2b2186aca2551aaa73b570bed35c043b;
key =      128'hafb394369ee4f0e24915324fa94e82fd;


#10;
 state = 128'hb2d470084854298ad5bc0a9a44a8180e;
key =      128'h8ef35bac9b2dd74c06e54209cdaf33c4;


#10;
 state = 128'h2d7f84a34776d4adec1c32def630c44a;
key =      128'h6c8523200407b2fbb90becf4c386ba20;


#10;
 state = 128'hecf1053eb73367d9e3a3509934d9d314;
key =      128'hf2a05ef705f6a810b4be0194fa7844bc;


#10;
 state = 128'h23e6694969da1ad07e4c7e6a48b32551;
key =      128'h943a5384909931fbee445732e5e9bc9b;


#10;
 state = 128'hf508cf25535ee2e9b2d2aa6054fa85d0;
key =      128'hd4e835d8986482667587a8d98a5a7065;


#10;
 state = 128'h2980623fa57cde4459574e89acad51d3;
key =      128'hec809586f185e417f1660c8cbb7cc07c;


#10;
 state = 128'h66e4fc22630b61da83bc62af3a2f69b4;
key =      128'h1627afff1f07ac9334116db84fef8d2d;


#10;
 state = 128'h63b6d489e4c7c135d8678324ec1296ed;
key =      128'hd80239459df80ae5a5d109771ff4c196;


#10;
 state = 128'hca82aa9590ae496cba6816cdf2a67aac;
key =      128'h99caa8b42a37c2b261cf08cb5e80c3c9;


#10;
 state = 128'hda28036e196ad74c99d3d2ed008b794c;
key =      128'hd49a5622e4fed118a345cdd9ff01c691;


#10;
 state = 128'h15d92ac9ee2f4301618702159e62137c;
key =      128'h8172fc69a66571cdcf49ab3e3ace4b71;


#10;
 state = 128'h764fa775ff647eeafd61eb81679bc3fe;
key =      128'h8ce90dbfbd324e7e6a8c7cf93ca45bc7;


#10;
 state = 128'hedb2f402f3ec167200f04d01cf678b10;
key =      128'h175b509998d48e9fd103610abe0da7bc;


#10;
 state = 128'h0eabbf9bd60198d5f6d6f2e516c53e7d;
key =      128'h2d2e218eb9c602af1f8ac9630cde9770;


#10;
 state = 128'h2b1a895607011b218bfdd80da4a1c216;
key =      128'h92d2cfe3354b98d2d155d561c2dd336c;


#10;
 state = 128'hdeedf7bc20e5ef13ddabe2c788814da4;
key =      128'hee1a531c4c2466eba81e793b686afbac;


#10;
 state = 128'h064658f30e262b47b2ebd20d3b3a6c1f;
key =      128'hab2a54c0f6f84eba739e16c704db0811;


#10;
 state = 128'ha70a22605bb5314d220da003cd5d470d;
key =      128'h5678879b9c4c70d5980fea86539cebf2;


#10;
 state = 128'h5afaa70ddbb5b0d85dfdc250a52a5a09;
key =      128'hb7fba3e29a544713233263315b76ce4e;


#10;
 state = 128'h4db6717571286b2137cf252e62dcf980;
key =      128'hb019d79c4f4a6d1e1f737cd1c07be94a;


#10;
 state = 128'h7b0d315acaed369cdb02bc5b523ddeb5;
key =      128'hd40257b695244cc412b597c8dbd23080;


#10;
 state = 128'hfd56e06171c84316b54dcaff5e078aa8;
key =      128'ha63309e11d3b57556e2ff0ee81490220;


#10;
 state = 128'hf87fa0e2e36947e3b998b61122189f41;
key =      128'hfdc84ba8901a04a215fe49f42d96484b;


#10;
 state = 128'hcb2515e86dae8f5c862746458da93fe5;
key =      128'h2c8a718a6abca475397fbaeeea671502;


#10;
 state = 128'h87b68c2b61f5641b90e71cabe51e905b;
key =      128'h7711a8023be1cd4d8a746087a174db76;


#10;
 state = 128'h83282a683ae41d8f94cacc395e79e85c;
key =      128'hded68a91df19b7578e698d18d12fdd69;


#10;
 state = 128'h97545708aed1397561439b0515c0bc84;
key =      128'h9ef39647657d0c4d02f3e699ccd322c4;


#10;
 state = 128'hef63287a669d346153c7e0cfe468879d;
key =      128'h6b825b1d01d00067aa03c4e66076d7e6;


#10;
 state = 128'h604fd9ffddc6ed0d6a308dcd324e9915;
key =      128'h5c9dd1f4b75d6ed1186260323679d837;


#10;
 state = 128'hbf96c8b2839c5cb5ffedcdea5a313c66;
key =      128'hdeb6cf0d6f95133dab87f77482e200d0;


#10;
 state = 128'h7e4178c9bf01ded511beefab386bef2b;
key =      128'hfb1622bea96aab357355f2a3bbf537f2;


#10;
 state = 128'h843a36afbf433b1455d0012aaf8d3cf1;
key =      128'h93aba35ef23d154ffa65920778b55ac9;


#10;
 state = 128'ha5fdef905564402b33ab3542cfe23871;
key =      128'h2b628ddcaa1d9fa3faa482316c735adc;


#10;
 state = 128'h74117049f2ca76b01c2575ab89eb08ad;
key =      128'h38b44d951ee3d1ed2f1987532b9c8ce1;


#10;
 state = 128'hac9fadfcce9f69238ceac4de6215d5cc;
key =      128'h109aca23ef2e7d9be61e4705cf11bad3;


#10;
 state = 128'h8b7cb168f95a1b1aac8544df3d0e9a1a;
key =      128'h004da8642bef7b2696110dc3306623c8;


#10;
 state = 128'heebbe2d4dce715fd74886c5a6bb19607;
key =      128'h656bfe3f3c905a7930d3a168986039c4;


#10;
 state = 128'h18871b1b8bf46e31e2ff7ddb524db013;
key =      128'h27b7b9ae7b644713adab37e98b460b70;


#10;
 state = 128'h58a3cd2716e3973b28f8e214407a4692;
key =      128'h126732ff628ecb79721039026cfd5645;


#10;
 state = 128'h5ec4a0234c75a7381b746d89b25befb3;
key =      128'h9ac5c22190fd538ed1030d8c863d0063;


#10;
 state = 128'hd9e401a1312559a87a4c9ac7aa2da789;
key =      128'hf844f26ad1884145b1a38b4e2d37e08c;


#10;
 state = 128'h8a061ce23cbc2b754eb708c51af8e4b0;
key =      128'h1b123dd6cdec9a7eb27e8f2652dfb670;

#10;
 state = 128'h7369c667ec4aff51abbacd2946e3fbf2;
key =      128'hf854c27c8de7e81b632e5a769ac99f33;


#10;
 state = 128'hb70d32665aa3583117055d25d45ee958;
key =      128'hc6cdb2ab1154b49b4174820e87dc3d21;


#10;
 state = 128'ha13ee97067fce141977e013e966bdcea;
key =      128'h2a5c388ffb3bb0ec543caf325cdb18ec;


#10;
 state = 128'h43fe1a023aaafafbe6d129fb947c3c05;
key =      128'h61bed875bb5cf989950f99a8b3f1ebb1;


#10;
 state = 128'h00f7ef05e53aa1e9d0cb0bcabd644748;
key =      128'ha81e231fc5647b1cc55a731463794b5e;


#10;
 state = 128'h2464703bdc099e11f2acd4aa3baf101b;
key =      128'h50e3cd335c15474819226fbbf57d9bba;


#10;
 state = 128'h1c1ae10b29f8237f131ba4f8e84ecab5;
key =      128'he0383298343d4d79774e5fbc056ccbfa;


#10;
 state = 128'h2b2186aca2551aaa73b570bed35c043b;
key =      128'hafb394369ee4f0e24915324fa94e82fd;


#10;
 state = 128'hb2d470084854298ad5bc0a9a44a8180e;
key =      128'h8ef35bac9b2dd74c06e54209cdaf33c4;


#10;
 state = 128'h2d7f84a34776d4adec1c32def630c44a;
key =      128'h6c8523200407b2fbb90becf4c386ba20;


#10;
 state = 128'hecf1053eb73367d9e3a3509934d9d314;
key =      128'hf2a05ef705f6a810b4be0194fa7844bc;


#10;
 state = 128'h23e6694969da1ad07e4c7e6a48b32551;
key =      128'h943a5384909931fbee445732e5e9bc9b;


#10;
 state = 128'hf508cf25535ee2e9b2d2aa6054fa85d0;
key =      128'hd4e835d8986482667587a8d98a5a7065;


#10;
 state = 128'h2980623fa57cde4459574e89acad51d3;
key =      128'hec809586f185e417f1660c8cbb7cc07c;


#10;
 state = 128'h66e4fc22630b61da83bc62af3a2f69b4;
key =      128'h1627afff1f07ac9334116db84fef8d2d;


#10;
 state = 128'h63b6d489e4c7c135d8678324ec1296ed;
key =      128'hd80239459df80ae5a5d109771ff4c196;


#10;
 state = 128'hca82aa9590ae496cba6816cdf2a67aac;
key =      128'h99caa8b42a37c2b261cf08cb5e80c3c9;


#10;
 state = 128'hda28036e196ad74c99d3d2ed008b794c;
key =      128'hd49a5622e4fed118a345cdd9ff01c691;


#10;
 state = 128'h15d92ac9ee2f4301618702159e62137c;
key =      128'h8172fc69a66571cdcf49ab3e3ace4b71;


#10;
 state = 128'h764fa775ff647eeafd61eb81679bc3fe;
key =      128'h8ce90dbfbd324e7e6a8c7cf93ca45bc7;


#10;
 state = 128'hedb2f402f3ec167200f04d01cf678b10;
key =      128'h175b509998d48e9fd103610abe0da7bc;


#10;
 state = 128'h0eabbf9bd60198d5f6d6f2e516c53e7d;
key =      128'h2d2e218eb9c602af1f8ac9630cde9770;


#10;
 state = 128'h2b1a895607011b218bfdd80da4a1c216;
key =      128'h92d2cfe3354b98d2d155d561c2dd336c;


#10;
 state = 128'hdeedf7bc20e5ef13ddabe2c788814da4;
key =      128'hee1a531c4c2466eba81e793b686afbac;


#10;
 state = 128'h064658f30e262b47b2ebd20d3b3a6c1f;
key =      128'hab2a54c0f6f84eba739e16c704db0811;


#10;
 state = 128'ha70a22605bb5314d220da003cd5d470d;
key =      128'h5678879b9c4c70d5980fea86539cebf2;


#10;
 state = 128'h5afaa70ddbb5b0d85dfdc250a52a5a09;
key =      128'hb7fba3e29a544713233263315b76ce4e;


#10;
 state = 128'h4db6717571286b2137cf252e62dcf980;
key =      128'hb019d79c4f4a6d1e1f737cd1c07be94a;


#10;
 state = 128'h7b0d315acaed369cdb02bc5b523ddeb5;
key =      128'hd40257b695244cc412b597c8dbd23080;


#10;
 state = 128'hfd56e06171c84316b54dcaff5e078aa8;
key =      128'ha63309e11d3b57556e2ff0ee81490220;


#10;
 state = 128'hf87fa0e2e36947e3b998b61122189f41;
key =      128'hfdc84ba8901a04a215fe49f42d96484b;


#10;
 state = 128'hcb2515e86dae8f5c862746458da93fe5;
key =      128'h2c8a718a6abca475397fbaeeea671502;


#10;
 state = 128'h87b68c2b61f5641b90e71cabe51e905b;
key =      128'h7711a8023be1cd4d8a746087a174db76;


#10;
 state = 128'h83282a683ae41d8f94cacc395e79e85c;
key =      128'hded68a91df19b7578e698d18d12fdd69;


#10;
 state = 128'h97545708aed1397561439b0515c0bc84;
key =      128'h9ef39647657d0c4d02f3e699ccd322c4;


#10;
 state = 128'hef63287a669d346153c7e0cfe468879d;
key =      128'h6b825b1d01d00067aa03c4e66076d7e6;


#10;
 state = 128'h604fd9ffddc6ed0d6a308dcd324e9915;
key =      128'h5c9dd1f4b75d6ed1186260323679d837;


#10;
 state = 128'hbf96c8b2839c5cb5ffedcdea5a313c66;
key =      128'hdeb6cf0d6f95133dab87f77482e200d0;


#10;
 state = 128'h7e4178c9bf01ded511beefab386bef2b;
key =      128'hfb1622bea96aab357355f2a3bbf537f2;


#10;
 state = 128'h843a36afbf433b1455d0012aaf8d3cf1;
key =      128'h93aba35ef23d154ffa65920778b55ac9;


#10;
 state = 128'ha5fdef905564402b33ab3542cfe23871;
key =      128'h2b628ddcaa1d9fa3faa482316c735adc;


#10;
 state = 128'h74117049f2ca76b01c2575ab89eb08ad;
key =      128'h38b44d951ee3d1ed2f1987532b9c8ce1;


#10;
 state = 128'hac9fadfcce9f69238ceac4de6215d5cc;
key =      128'h109aca23ef2e7d9be61e4705cf11bad3;


#10;
 state = 128'h8b7cb168f95a1b1aac8544df3d0e9a1a;
key =      128'h004da8642bef7b2696110dc3306623c8;


#10;
 state = 128'heebbe2d4dce715fd74886c5a6bb19607;
key =      128'h656bfe3f3c905a7930d3a168986039c4;


#10;
 state = 128'h18871b1b8bf46e31e2ff7ddb524db013;
key =      128'h27b7b9ae7b644713adab37e98b460b70;


#10;
 state = 128'h58a3cd2716e3973b28f8e214407a4692;
key =      128'h126732ff628ecb79721039026cfd5645;


#10;
 state = 128'h5ec4a0234c75a7381b746d89b25befb3;
key =      128'h9ac5c22190fd538ed1030d8c863d0063;


#10;
 state = 128'hd9e401a1312559a87a4c9ac7aa2da789;
key =      128'hf844f26ad1884145b1a38b4e2d37e08c;


#10;
 state = 128'h8a061ce23cbc2b754eb708c51af8e4b0;
key =      128'h1b123dd6cdec9a7eb27e8f2652dfb670;


#10;
 state = 128'h47dce5d2d684981051243ba1f56b1d1f;
key =      128'hd8107d5a3da5fc17fcef248cac4eceda;


#10;
 state = 128'hc4f32ab3649a77c3d1b5beb235c620db;
key =      128'hb40ed69d5ff2b3d3b15be1d7635da9b0;


#10;
 state = 128'h962751d37bfac1c85b4caf806c9113cf;
key =      128'hbc219fe92a1b1352a4db76f4f308391f;


#10;
 state = 128'h52892f8a71cd84f103cc1a33166f5d2d;
key =      128'h4fd390fc9879eea3843c54651777448d;


#10;
 state = 128'h656a0174b8d637857ebba251fc952b00;
key =      128'h5f4b68bbbbf7c456a6403319ecbeb778;


#10;
 state = 128'h3d5128b8b1f6275fc92fb1c998c6c4dc;
key =      128'h83f7112cef3eeed699957e21ee855336;


#10;
 state = 128'hdb2cd67bc78c22fdb090bbd3ac485680;
key =      128'h3e2f3f684e2d6e2d22e8c2ec91116d16;


#10;
 state = 128'h416c3d443208f85f34e299b457e02aef;
key =      128'h969510696ae5c27e9b8dcd857e2c9e3a;


#10;
 state = 128'h3ac099db456cc89151794f61e3a85a79;
key =      128'he8793e6a85525e006620df2b58e44d7d;


#10;
 state = 128'h7792a4e6cebdff6dc71f364efaaac890;
key =      128'h06e22406ae8c35829214ac14dfeaf8f9;


#10;
 state = 128'h0a577d9dcad8147cdb91f84ac6d53cc0;
key =      128'he2ccb860019058edfe93a4053ade7e9d;


#10;
 state = 128'h774435fb93411c49d46ed2146e9a440e;
key =      128'he95167fcc4eae1bf23c37e86f75da1fc;


#10;
 state = 128'h1f6ea1d6d2b2afbd90a6218161fe4165;
key =      128'h674a4fa8b72c3431aedaefb266a53790;


#10;
 state = 128'h958513d8446737c2bdd40e58f71ed24f;
key =      128'h535e68224f0a8a9d09fee479f36fa31b;


#10;
 state = 128'h7988f4b784bdf02c4d4291fe86446064;
key =      128'h66d9a2c9a6b5e32de2b0b3c70ed51f57;


#10;
 state = 128'h40875d144bc4454d3a9806d630c0dc67;
key =      128'hac96997f43524b7c562502ff3664fa22;


#10;
 state = 128'ha576eb5807f13a30a8418941e5d80266;
key =      128'h18916e9bb85be3b9080e81e6d33e727b;


#10;
 state = 128'h8e79b45e2f956aee59d7d7f3743eafd9;
key =      128'hd78ccf1d998fe8b3e4a19e696eb8df10;


#10;
 state = 128'h81fd31938eb1929b42e8886955b72638;
key =      128'ha92c43f69442bc2b6a79e35a55d931c2;


#10;
 state = 128'hfdd6d662d28b876848147310909dcb9a;
key =      128'h3a39ca0fe0cf7b86204a485edb752379;


#10;
 state = 128'h62d84bf9e33463d3712b48d72301c814;
key =      128'h185d3a9213f82cb5ed33437460c8a866;


#10;
 state = 128'hc6c2a0f3dba9f604524cd43e2f754d9d;
key =      128'h3c48d387744f40ffea6182831d4a2a2a;


#10;
 state = 128'hcee40cca40a98d02ff93f562c92e0842;
key =      128'hdb0576db3a4f54b70024b0d6a51e6eda;


#10;
 state = 128'h7c73027af1bd1d8f55f05012341e1f58;
key =      128'h4c0f24954f875e78e94fab0e948e6d1a;


#10;
 state = 128'hff11016f31f0ce1e7686e11e95aaa400;
key =      128'h41e2b9c8269069172e0fdf14bcc39d4d;


#10;
 state = 128'hbdbbd49ec0eeaca28d36748de122e118;
key =      128'hb222049a82d8b26ddeb0e791229b7384;


#10;
 state = 128'he9df56478fa9cd025a1ce0415b3b3fc1;
key =      128'hb10d5d43a033e50f507fe3cc9e731a57;


#10;
 state = 128'h7388527061023120d2bb1f11a12ef65e;
key =      128'h62523b53ed038521c03e82690c5eb19c;


#10;
 state = 128'h237fe60329858218fffc40a18aa02a37;
key =      128'h86edf365e174f0780ea1b272661a0063;


#10;
 state = 128'hfe8a9ae6bd280f1c86bc244fb3115c4e;
key =      128'hc83afe4f60a9aeeec36e4b603129884b;


#10;
 state = 128'h3e30b32212fb58c2ca98b77c637da914;
key =      128'h952bb7a7c5f5d5656b8863200e9cb2ec;


#10;
 state = 128'h284dcc65a03a4824146ad2002377e87c;
key =      128'h05b9a39f98caae78fe0353126a0c9f05;


#10;
 state = 128'h9092596ca231cca21bb69b9f233e2d83;
key =      128'h4828f7d0b8e0f2a64ab6e345efb5c283;


#10;
 state = 128'hbe7f471cb360b014cfce164c14f20c43;
key =      128'haa5c1a0452623d0da39d1820f69252da;


#10;
 state = 128'hadb412990e6014c26ede2e2a3f82d03b;
key =      128'hf8e9deeb3c4a4b1b3ddfe763d3347239;


#10;
 state = 128'h4680e8842755e1fd4a95330fee891703;
key =      128'h11e672f6204d31bd525e2d182325929f;


#10;
 state = 128'h7769a57a969fbe86f5e034f142e36a4c;
key =      128'h9a53cadc13baa1fb6d6518ce25908aaa;


#10;
 state = 128'hb69cf930a94c3bb8bc9e2d7073fe8297;
key =      128'h470d514cc05ac8f28b2dc0e07ab0bd4a;


#10;
 state = 128'h6f314cb7f8187d8841b4b7aa85b5b239;
key =      128'hf6ccc2036bb6268a31f6e4e658aba6a1;


#10;
 state = 128'h7ac7dcf20472e05ad0462697dc55fbd8;
key =      128'h48d221bd2eb388470e5fa96c41660a4f;


#10;
 state = 128'h41bc2ee7a5452e0e2d758b554409ca86;
key =      128'h328cdbebd0603f6437debfe8b17845ca;


#10;
 state = 128'h81f23473b826376349e59bc3508def65;
key =      128'h2e8219ca40ffe3586c77dda2951df022;


#10;
 state = 128'h87160f240a3f3c473c5325d7de8ce114;
key =      128'h530d0ffa94930cf20c010be91fa11efb;


#10;
 state = 128'h75a7b82ecc7fe6f41f08d20baefe95b3;
key =      128'h96010ba4002a94179a0c2b9f78baae4a;


#10;
 state = 128'h5aed616653266c47f2722f3e68a070c4;
key =      128'h92fea17bd59328359e6f9f54b316294d;


#10;
 state = 128'hd20e038aad25346f279f9763838f3f08;
key =      128'h16168de00aeba9b696a85a480e49be84;


#10;
 state = 128'h30e057c1efdd058ca5177d9d9d28a6bc;
key =      128'heab33e3430f49ee77cc69cf81b8b0f5a;


#10;
 state = 128'hf34b6b670ee2287162b3f9a5d4ffdba0;
key =      128'h01beb21a4831b250a8c5f74e6ec35007;


#10;
 state = 128'h2c610ebbdc3a4336dd3eed3de3b13dc9;
key =      128'h3fe46fef6f87162114174c0d5882da9c;


#10;
 state = 128'h1e84e3e864fabf27754138ac6458f275;
key =      128'h82a33d6160f12b5314750877ca6cf7e2;


#10;
 state = 128'h02e8f0db5c66e3af91d1a71bfaf52a99;
key =      128'hba7c99673b1a6dc4574f8f756221bb87;


#10;
 state = 128'h5b6409ac08b7caec0a9989711a048eb3;
key =      128'hebd480276227eeed05b9767ede67da32;


#10;
 state = 128'hd039cbe306d8f1952d10717a274714ff;
key =      128'h81121b9487e33909e28c9cb059c0f376;


#10;
 state = 128'h5329f9be645901ea729169721199d87d;
key =      128'hfd92abf3958475e587771111c3e13704;


#10;
 state = 128'h1b160a307e7f700c57f011d9dd6889e9;
key =      128'h1adafb3582af5e707409266f8d37ea5d;


#10;
 state = 128'h01a84df5977f28bd22ee70392eff56f9;
key =      128'hc248d951a744f7387a1b4d1d2d085238;


#10;
 state = 128'h5d2eb0a011f4add81734e21d8a453339;
key =      128'h454c8e0da3ec9085161d08defa43255a;


#10;
 state = 128'hae5871d63cc04c1e6853f42f34f29827;
key =      128'hac793f26ad4f66cfc8c36c6e68c30692;


#10;
 state = 128'h96161b7796d2d667f2fe25cae426f1bd;
key =      128'hff90a03074addf06dd3c704bee45ff77;


#10;
 state = 128'h82845c1afd18563239ef177b381d1508;
key =      128'hbb37adb5d72fe48cccb56c5586bafa6b;


#10;
 state = 128'h89083f56118620953f4a75374077678a;
key =      128'ha0fbaf14e8772b9302b42c977d886f27;


#10;
 state = 128'h430690aee8548cb18c289e0119cc9f05;
key =      128'he2b9c74e89ca31f2848c7f5d9c0214ee;


#10;
 state = 128'h56df08a5963e3495d82266d254f1ee06;
key =      128'ha836abb6393201dc6ebebe80770ac0d2;


#10;
 state = 128'h5dcde9c8f0f40c1d78c81672bbcdb905;
key =      128'h40630364847a950426f23853c09dfcf8;


#10;
 state = 128'h031e6be6e9f312772d62bb28d9e82f75;
key =      128'h371a4c3235bb94e1c45baecc9084f8aa;


#10;
 state = 128'hda94a263ddc487b4b80a26438791f355;
key =      128'h20beab3f0b557a3fd2cfb0280c6354a9;


#10;
 state = 128'habe7f7f6c188ab7e267992d1c4ad0b85;
key =      128'hf6e56cb60e013ae694e0d1eb1ba04325;


#10;
 state = 128'hb9c6873a037a4e326629f4e1b52bd7ff;
key =      128'h29ab10433537ad4aa3c9177e95be6a5b;


#10;
 state = 128'h244e85f1b427c9d3bc1b51bd6b714628;
key =      128'ha0941d5648d6cbca3deb9fe2fbd3a909;


#10;
 state = 128'h021f212ea7b646eabf63d1976d2ad517;
key =      128'hbc0ebef26c04e4898da9ef83c7887c98;


#10;
 state = 128'h88c9a79e85307fed684493515ad66f68;
key =      128'hb716e42d4b231ac8a2d8cc09e7696049;


#10;
 state = 128'hf56f3207027a9fb19b6bbe335bf6412d;
key =      128'hed120c25303835274ad2110179313b71;


#10;
 state = 128'h1f6ea16d7321e840d40f8ca6f22f05cd;
key =      128'h38df4111776918769ac23b29e413f377;


#10;
 state = 128'hd5038194104825697fe457b16e71135c;
key =      128'hcaa6515492410f69c22c034b8ba640f7;


#10;
 state = 128'h2b60aac1803ba9cf5dff1f0086cb7132;
key =      128'h2b5071c2ccbd91818c8ee995eb173429;


#10;
 state = 128'had1678de212e5121a27e2d706028499e;
key =      128'h3c8b78bb9e0848095b2a9632a94642ca;


#10;
 state = 128'hdb565cba1dfc84ad50bf7bb27fb1e7c4;
key =      128'h69bb3c5fb707c385241232592ecd5974;


#10;
 state = 128'h630923b55a8005a845aa408087c45b27;
key =      128'h1df080989dd4f7439dc1e629f5cb8e3f;


#10;
 state = 128'h5958d4b15ab3d8da409f5e1851c764b9;
key =      128'h276eb7e4d8c442ae68758529c55d4113;


#10;
 state = 128'hef1eb515a64ad28ee9e6e930313bad4d;
key =      128'h1359a96415eb1decb67d60a3b77bdba1;


#10;
 state = 128'h1ea69a909cc5f06c2785abdabd59c059;
key =      128'h56d0b26a726bbbcfbd29e81c5474a4c3;


#10;
 state = 128'haa721b3ee546370b3c0dcce3f6f9668c;
key =      128'he74cca18a15ab785635f83a066b7d327;


#10;
 state = 128'hfa102aee44df5761af80ec236aa67a52;
key =      128'hc952f2444a6bacaa56adca2f8cbc659d;


#10;
 state = 128'hf086cd8f47356524a4f6b552730f9c2f;
key =      128'h393d618f3c83a80d0f923072249b4f95;


#10;
 state = 128'h4015211cd9874a872f7d7dffa9a28c1a;
key =      128'hfae2dfedf93665872b09c995344fa418;


#10;
 state = 128'h4d7464c6ae26fbae92dda3781d3b7f30;
key =      128'he6181d5f18e04e822f43e9175363928d;


#10;
 state = 128'ha5a0d7f74b53c6d29add306a0fb719b0;
key =      128'hb9f5cf3635d1d51e4c6514be9d9fc8a6;


#10;
 state = 128'h724340a070bd9606770a9bc7ea86c2b4;
key =      128'hafa37b910fe574512f5b4a88b2ccfb12;


#10;
 state = 128'h41250f3b6db2e2a631e4bc7d101c6a7e;
key =      128'h36bfbfe5bc46a43401eba1eed7b3b89c;


#10;
 state = 128'h6d19d8c738dacbbb066abe870e168628;
key =      128'h7944d54568368a7ac869212ca1a01dd9;


#10;
 state = 128'hb00eb9f50be9e984d01153a71ede27d9;
key =      128'h779822fdd9dfceadc9a149ef5b6a4166;


#10;
 state = 128'h7e0c78fa098af56121d99b48c03fb7c3;
key =      128'h8637d7d9955f16a5c55e015f3d21c842;


#10;
 state = 128'ha2bb2d406aab4522a48b84e11464ca3b;
key =      128'h479b9ba211dcfab13ed63afb437bf702;


#10;
 state = 128'h46e536245db0907c4f013b14a8636506;
key =      128'hb1effe00f4c2ccf909329906b54cad90;


#10;
 state = 128'h60fb31e4d5bdacc1ed24bee723958723;
key =      128'h7fd4858657739751c060a6303775ac53;


#10;
 state = 128'h9e9771dd0473541d35f29712a558871f;
key =      128'h5d242d0cf4b597c491b4153d9fc82ac2;


#10;
 state = 128'hb83e609bc7bcb1b468fcae49420d5536;
key =      128'h46a03182063a55c82c97ee6ab3cc5f18;


#10;
 state = 128'h746b0abf043b28bb0c6c37d60e4f798c;
key =      128'h7354efaaae798e4495db107d2f49a76f;


#10;
 state = 128'h6ca3b4b1b371dedca2bfdd1501b00e57;
key =      128'h417405fd10f0ed936da6cbfd239cef72;


#10;
 state = 128'h808f3fa33233001d35d4f2defe368501;
key =      128'h1d40ab8a962e30986d03d4fb66909fc3;


#10;
 state = 128'hfbe61fdefe2d19200d33020c110b6987;
key =      128'had2e4b1476435c7bf3e34630c35a73e5;


#10;
 state = 128'hb3be409366b1eb5a7473e4ed62857e4d;
key =      128'h450fb4ca41bc52107d349f98a6408e13;


#10;
 state = 128'h2959fecfd78f0ae93b4b02ee4a9dd180;
key =      128'h9590ac8596d64cfefe130beb68a45399;


#10;
 state = 128'h3b91fd51f5122007a3315d22b3edce2e;
key =      128'h79497d7bb5101fc9c4b3232ac82c5877;


#10;
 state = 128'h5d03be55015215dea1a48373cd559152;
key =      128'hd8469e0fe88d56bdf1ac417aeeb9d899;


#10;
 state = 128'h754bbd9645769ed273e71a21ba403cab;
key =      128'h979387da577f20ddfa482b619ae90204;


#10;
 state = 128'h910f34bff4d785d24b67be9fd405a8fa;
key =      128'h0c6b982f1a64ebb91a15ac166db5feae;


#10;
 state = 128'h05ffc432e9f9d64a8e34609437623a08;
key =      128'h8b44cdd2cfa6a8b803e9bb54eb709eb9;


#10;
 state = 128'hadf06f63d996e9455267cb4ad78ac905;
key =      128'h4f63ce97ca1e09767dcd08c409683ea6;


#10;
 state = 128'hf3b659ad8ccc4d421ddf341894f469fd;
key =      128'hade4573724770260b1a1450a30ba0a83;


#10;
 state = 128'ha5237163d632f0be21f31124b1b6e77a;
key =      128'h9f5e9a3fa7c4d59c9d58651ad2ce126f;


#10;
 state = 128'h4178f1830517aae135270abb31e6ddf2;
key =      128'h13d0447734ba941969d112faa83c9f25;


#10;
 state = 128'h72eab4911978015efe4e9f0cf32f347c;
key =      128'h9106ff788ec5c194f8f797d3c7a13336;


#10;
 state = 128'h453a8be7985eb28ccd96ac5158c0c5e0;
key =      128'h59eac6c55be7af877d53de46f944f412;


#10;
 state = 128'h0c3f7e7f81a49d302a4e3b4ac5830e00;
key =      128'h5c1e6dd563b7051cf6e00be47fef24ff;


#10;
 state = 128'hd38b2ea316552fcc6b40a36a8730c3b2;
key =      128'h4de34f3038b09b54a52e90a657241eb4;


#10;
 state = 128'h182baf4c492e80dfd5b46f23635ce532;
key =      128'h88b0403481c160dba426eff05afc4b0d;


#10;
 state = 128'hd97227faca23a1a742a0d710f0a5fcbc;
key =      128'h1779553ca5983ab5374abf290491460a;


#10;
 state = 128'h14de036db4de01a495f77ed8b7859c7b;
key =      128'ha7cffef2624d6738309997264a352add;


#10;
 state = 128'hd25e132dec863c1436817dbb0ced071a;
key =      128'h3eb3bc054aa00024747b399790beb063;


#10;
 state = 128'hd7621cc314c3e959804a4566518c374c;
key =      128'h188f40f4d8622f40cb4cdd68505c0b8d;


#10;
 state = 128'h8027be270e94eba77c8ede300acd1b16;
key =      128'h9b225d5bf573848cefc0c062f2401ccb;


#10;
 state = 128'h827367db82900752fcfe1fe69506cc3a;
key =      128'hb53028290eaaa4ac2ffe6b6462213e87;


#10;
 state = 128'hf8e594a5827a759cce7e79946e638445;
key =      128'h582394ac9c67ce38c0cb65394823eca3;


#10;
 state = 128'h1d400881129fbb7d79e01d344de744a1;
key =      128'h10a50ad811ac0cd814d27771e45df563;


#10;
 state = 128'h7a019dfd8c8ca0585e056dbd89abecb1;
key =      128'hcf9951f7cfe1455d1fe3b3bca50440a8;


#10;
 state = 128'h361f05de63c3aca6cac2c819ac536db5;
key =      128'h1c7becbeedeb5c31b70cce0fed5c100f;


#10;
 state = 128'hbc237c16411fe628640be1af0d105e4f;
key =      128'h7b298b4af76814e8f2af74e39bdf0b85;


#10;
 state = 128'haf57028798f076e9a7fcfb58a3b40c59;
key =      128'h7f1ede97d57786f280c726fbb91ba631;


#10;
 state = 128'h926872a9402a59e8aee72654c9519c32;
key =      128'h6c49707af142c0f6177109e659d08cb0;


#10;
 state = 128'he7eb39fee62715926d940f3b2536e6ab;
key =      128'h4c917f56253ed33f8d3dafdd3ae60d3c;


#10;
 state = 128'hd821d14621bf49e6038e53588f28c439;
key =      128'h83dcb9446aa91a8d05f7e6c93a40ddf3;


#10;
 state = 128'h941261ae02b5d1aa5e0543254bee2d07;
key =      128'h74cfcae7adde78e451b3d55e608bf3b2;


#10;
 state = 128'hfff49e549401a96ff3f307ec1b3fe134;
key =      128'h8f8f0eabe43c6d86f435ef423754c1e2;


#10;
 state = 128'hce36485fdd6337f173d1563ee28e1037;
key =      128'ha4711e1ece88ad8b7fc2bd9dddb6177e;


#10;
 state = 128'h51acec5f622e0f249cd5ff652d7e640f;
key =      128'h0dd1ef8239db599c95b99e1714736fb5;


#10;
 state = 128'h80651f5c93e2942ea32fb8939ed0ad1c;
key =      128'h38aba29c127287fbdaa82b25f6ee1b9a;


#10;
 state = 128'h6876543a7bfb59e82d1e2a1173cbefd7;
key =      128'h8cab7691229f1dfde3fc47489cd9eb62;


#10;
 state = 128'h2704503fbaa2ffa900e7c1294173b2b0;
key =      128'h26cd1e2884486c3c156745b36fb14130;


#10;
 state = 128'h3a96b591ddf438b4a9dddbf9b5ea508d;
key =      128'habdbb86fd82f242499ed976969089fd8;


#10;
 state = 128'h09a39e54d0e697d6ff79c47283b46414;
key =      128'h402e901c1d185eb4cdb606f5f936bea5;


#10;
 state = 128'h3202d95ce202e970c1e17cadfc4595e0;
key =      128'hd93c7325c6f655d10093ac5bc6f9c96a;


#10;
 state = 128'h12f9fca292f4fbe55753d5779053986b;
key =      128'hdd6a900c40a460e57740370da33e3901;


#10;
 state = 128'h1ab63735aaacaa32eb010080a47b5598;
key =      128'hca82e5e5530a26465eca4a5db9020883;


#10;
 state = 128'h72d3b83fe21c806218cd1d8057bd4972;
key =      128'h74213f2ec2c72b65f9219275dab2239a;


#10;
 state = 128'h3d4c85db85206805f89eed85654f5b36;
key =      128'hffd9719a12c1a19ccd0be233e0a7bd05;


#10;
 state = 128'h481ef342e1cd3e5b62d96b2b60c728c6;
key =      128'h365fa099744821410942530352e9e910;


#10;
 state = 128'h389a07dd711968459ad3f2d3b4fa9a1b;
key =      128'h7cea5a3a7ef0327b95873285f9e8711c;


#10;
 state = 128'hbe318278be2f4bea5858023dd60d529c;
key =      128'h2752f7acafa6432a91452d75178a2d9e;


#10;
state = 128'h9ad5bcaf44580407a29db006af78aa02;
key =      128'hcbd6cba1837b7c0e4815c0aa9c5f9fed;
#170;

$display("Good.");
//
#100
$finish;
end
  
  initial begin 
    $dumpvars;
    $dumpfile("waves_aes_128.vcd");
  end
    always #5 clk = ~clk;
endmodule

